vhdl/Week1/AAC2M1P1/aac2m1p1_types.vhdl