vhdl/Week1/AAC2M1P1/AAC2M1P1.vhdl